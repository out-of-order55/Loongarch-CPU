module bjp_unit(
    
);

endmodule